    Mac OS X            	   2   �      �                                      ATTR       �   �   #                  �   #  com.apple.quarantine q/0082;5d6f0d88;The\x20Unarchiver; 